// code converter

module code_conv_7seg
(
input [3:0] x,
output reg [0:7] y
);

always @(x)
begin 
	case(x)
		4'b0000: y=8'b00000010;
		4'b0001: y=8'b10011110;
		4'b0010: y=8'b00100100;
		4'b0011: y=8'b00001100;
		4'b0100: y=8'b10011000;
		4'b0101: y=8'b01001000;
		4'b0110: y=8'b01000000;
		4'b0111: y=8'b00011110;
		4'b1000: y=8'b00000000;
		4'b1001: y=8'b00011000;
		4'b1010: y=8'b00010000;
		4'b1011: y=8'b00000000;
		4'b1100: y=8'b01100100;
		4'b1101: y=8'b01100000;
		4'b1110: y=8'b00000010;
		4'b1111: y=8'b01110000;
		default: y=8'bx;
	endcase
end
endmodule
